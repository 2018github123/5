// testbench_top:
//              This is the top most file,which connects the DUT and TestBench
//              TestBench top consists of DUT,Test and Interface instance
//              Interface connects the DUT and TestBench

module testbench_top;

bit clk;
bit reset;


endmodule