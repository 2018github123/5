`timescale 1 ns / 100 ps
