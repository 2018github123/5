program env(intf.env if1);
    clocking cb @(posedge if1.clk);
        output select = if1.select;
        input dtoe = if1.dtoe;
        output etod = if1.etod;
        inout bus = if1.bus; 
    endclocking
    
    covergroup cov @cb;
        //slt_cp:coverpoint cb.select;
        dte_cp:coverpoint cb.dtoe;
        //etd_cp:coverpoint cb.etod;
        bs_cp:coverpoint cb.bus;
        cs_cp: cross dte_cp,bs_cp;
        option.per_instance = 1;
    endgroup

    task doit(input logic [1:2] sel, input logic [1:4] toe,bd);
        cb.select <= sel;
        cb.etod <= toe;
        cb.bus <= bd;
    endtask

     initial begin
        cb.etod <= 4'b0000;
        cb.bus <= 4'bz;
        @cb doit(2'b00, 4'b1001, 4'bzzzz);
        @cb doit(2'b01, 4'b0110, 4'bzzzz);
        @cb doit(2'b10, 4'b0101, 4'b01x1);
        @cb doit(2'b11, 4'b0001, 4'bzzzz);
       // @cb $finish(0);
      end

      initial forever @cb begin
        $display("at %0d, in %m: select=%b etod=%b dtoe=%b bus=%b", 
          $time, if1.select, if1.etod, if1.dtoe, if1.bus);      
      end
      
     initial begin 
        cov cg = new();
        if(cg.dte_cp.get_inst_coverage <= 33.33)
         begin
            $write("cov = %3.5f \n",cg.dte_cp.get_inst_coverage());
         end
     end
endprogram
